// ##############################################################################
// ## Intel Top Secret                                                         ##
// ##############################################################################
// ## Copyright (C) Intel Corporation.                                         ##
// ##                                                                          ##
// ## This is the property of Intel Corporation and may only be utilized       ##
// ## pursuant to a written Restricted Use Nondisclosure Agreement and any     ##
// ## applicable licenses with Intel Corporation.  It may not be used,         ##
// ## reproduced, or disclosed to others except in accordance with the terms   ##
// ## and conditions of such agreement.                                        ##
// ##                                                                          ##
// ## All products, processes, computer systems, dates, and figures            ##
// ## specified are preliminary based on current expectations, and are         ##
// ## subject to change without notice.                                        ##
// ##############################################################################
// ## Text_Tag % __Placeholder neutral1

module ctech_lib_clk_nand_en (
   input logic clk,
   input logic en,
   output logic clkout );

   logic 	clkout_and;
   g1iclb0a2ab1n04x5 ctech_lib_clk_nand_en_dcszo1 (.clk(clk),.en(en),.clkout(clkout_and));
   g1icinv00ab1n04x5 ctech_lib_clk_nand_en_dcszo (.clk(clkout_and), .clkout(clkout));

endmodule // ctech_lib_clk_nand_en
