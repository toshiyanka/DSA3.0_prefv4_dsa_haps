// ##############################################################################
// ## Intel Top Secret                                                         ##
// ##############################################################################
// ## Copyright (C) Intel Corporation.                                         ##
// ##                                                                          ##
// ## This is the property of Intel Corporation and may only be utilized       ##
// ## pursuant to a written Restricted Use Nondisclosure Agreement and any     ##
// ## applicable licenses with Intel Corporation.  It may not be used,         ##
// ## reproduced, or disclosed to others except in accordance with the terms   ##
// ## and conditions of such agreement.                                        ##
// ##                                                                          ##
// ## All products, processes, computer systems, dates, and figures            ##
// ## specified are preliminary based on current expectations, and are         ##
// ## subject to change without notice.                                        ##
// ##############################################################################
// ## Text_Tag % __Placeholder neutral1

module ctech_lib_clk_nor_en (
   input logic clk,
   input logic en,
   output logic clkout );

   logic clkout_or;
   g1iclb0o2ab1n04x5 ctech_lib_clk_nor_en_dcszo1 (.clk(clk),.enb(en),.clkout(clkout_or));
   g1icinv00ab1n04x5 ctech_lib_clk_nor_en_dcszo (.clk(clkout_or),.clkout(clkout));
   
endmodule // ctech_lib_clk_nor_en
